`ifndef TIMEALIGN_UVC_PKG_SV
`define TIMEALIGN_UVC_PKG_SV

package timeAlign_uvc_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;


  `include "timeAlign_uvc_agent.sv"

endpackage: timeAlign_uvc_pkg

`endif  //TIMEALIGN_UVC_PKG_SV